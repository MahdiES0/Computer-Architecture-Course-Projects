module MazeTb();
    
    MyMaze M1(start, clk, rst, run, fail, done, move);
endmodule